
entity VOTE_SELECTOR is
  port(
    head_ref: in std_logic;
    ref_1 : in std_logic;
    ref_2 : in std_logic;
    ref_2: in std_logic;
    vote: out std_logic

    );

end VOTE_SELECTOR

  signal 
archtecticture ARCH_VOTE_SELECTOR of VOTE_COUNTER is 
  begin
    
